IP_CORE_PLL_inst : IP_CORE_PLL PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
